library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity ROM_176x4 is
  port (--Clock : in std_logic;
  		CS_L : in std_logic;
        R_W  : in std_logic;
        Addr   : in std_logic_vector(7 downto 0);
        Data  : out std_logic_vector(3 downto 0));
end ROM_176x4;

architecture ROM_176x4_Arch of ROM_176x4 is
  type rom_type is array (0 to 175)
        of std_logic_vector (3 downto 0);
  signal ROM : rom_type;
  signal Read_Enable : std_logic;
begin

ROM(0) <= X"5";
ROM(1) <= X"0";
ROM(2) <= X"4";
ROM(3) <= X"2";
ROM(4) <= X"3";
ROM(5) <= X"D";
ROM(6) <= X"0";
ROM(7) <= X"B";
ROM(8) <= X"5";
ROM(9) <= X"1";
ROM(10) <= X"4";
ROM(11) <= X"3";
ROM(12) <= X"3";
ROM(13) <= X"D";
ROM(14) <= X"1";
ROM(15) <= X"B";
ROM(16) <= X"8";
ROM(17) <= X"0";
ROM(18) <= X"B";
ROM(19) <= X"D";
ROM(20) <= X"4";
ROM(21) <= X"B";
ROM(22) <= X"F";
ROM(23) <= X"0";
ROM(24) <= X"B";
ROM(25) <= X"3";
ROM(26) <= X"D";
ROM(27) <= X"0";
ROM(28) <= X"B";
ROM(29) <= X"F";
ROM(30) <= X"1";
ROM(31) <= X"B";
ROM(32) <= X"3";
ROM(33) <= X"D";
ROM(34) <= X"1";
ROM(35) <= X"B";
ROM(36) <= X"8";
ROM(37) <= X"0";
ROM(38) <= X"B";
ROM(39) <= X"D";
ROM(40) <= X"5";
ROM(41) <= X"B";
ROM(42) <= X"F";
ROM(43) <= X"0";
ROM(44) <= X"B";
ROM(45) <= X"C";
ROM(46) <= X"1";
ROM(47) <= X"B";
ROM(48) <= X"D";
ROM(49) <= X"8";
ROM(50) <= X"B";
ROM(51) <= X"F";
ROM(52) <= X"0";
ROM(53) <= X"B";
ROM(54) <= X"3";
ROM(55) <= X"D";
ROM(56) <= X"0";
ROM(57) <= X"B";
ROM(58) <= X"F";
ROM(59) <= X"1";
ROM(60) <= X"B";
ROM(61) <= X"3";
ROM(62) <= X"D";
ROM(63) <= X"1";
ROM(64) <= X"B";
ROM(65) <= X"8";
ROM(66) <= X"0";
ROM(67) <= X"B";
ROM(68) <= X"D";
ROM(69) <= X"6";
ROM(70) <= X"B";
ROM(71) <= X"F";
ROM(72) <= X"0";
ROM(73) <= X"B";
ROM(74) <= X"C";
ROM(75) <= X"1";
ROM(76) <= X"B";
ROM(77) <= X"D";
ROM(78) <= X"9";
ROM(79) <= X"B";
ROM(80) <= X"F";
ROM(81) <= X"0";
ROM(82) <= X"B";
ROM(83) <= X"3";
ROM(84) <= X"D";
ROM(85) <= X"0";
ROM(86) <= X"B";
ROM(87) <= X"F";
ROM(88) <= X"1";
ROM(89) <= X"B";
ROM(90) <= X"3";
ROM(91) <= X"D";
ROM(92) <= X"1";
ROM(93) <= X"B";
ROM(94) <= X"8";
ROM(95) <= X"0";
ROM(96) <= X"B";
ROM(97) <= X"D";
ROM(98) <= X"7";
ROM(99) <= X"B";
ROM(100) <= X"F";
ROM(101) <= X"0";
ROM(102) <= X"B";
ROM(103) <= X"C";
ROM(104) <= X"1";
ROM(105) <= X"B";
ROM(106) <= X"D";
ROM(107) <= X"A";
ROM(108) <= X"B";
ROM(109) <= X"F";
ROM(110) <= X"0";
ROM(111) <= X"B";
ROM(112) <= X"E";
ROM(113) <= X"1";
ROM(114) <= X"B";
ROM(115) <= X"4";
ROM(116) <= X"0";
ROM(117) <= X"F";
ROM(118) <= X"7";
ROM(119) <= X"B";
ROM(120) <= X"B";
ROM(121) <= X"9";
ROM(122) <= X"A";
ROM(123) <= X"F";
ROM(124) <= X"A";
ROM(125) <= X"B";
ROM(126) <= X"B";
ROM(127) <= X"4";
ROM(128) <= X"8";
ROM(129) <= X"9";
ROM(130) <= X"2";
ROM(131) <= X"A";
ROM(132) <= X"F";
ROM(133) <= X"6";
ROM(134) <= X"B";
ROM(135) <= X"B";
ROM(136) <= X"9";
ROM(137) <= X"A";
ROM(138) <= X"F";
ROM(139) <= X"9";
ROM(140) <= X"B";
ROM(141) <= X"B";
ROM(142) <= X"3";
ROM(143) <= X"9";
ROM(144) <= X"9";
ROM(145) <= X"2";
ROM(146) <= X"A";
ROM(147) <= X"F";
ROM(148) <= X"5";
ROM(149) <= X"B";
ROM(150) <= X"B";
ROM(151) <= X"9";
ROM(152) <= X"A";
ROM(153) <= X"F";
ROM(154) <= X"8";
ROM(155) <= X"B";
ROM(156) <= X"8";
ROM(157) <= X"4";
ROM(158) <= X"B";
ROM(159) <= X"B";
ROM(160) <= X"9";
ROM(161) <= X"A";
ROM(162) <= X"7";
ROM(163) <= X"0";
ROM(164) <= X"4";
ROM(165) <= X"1";
ROM(166) <= X"9";
ROM(167) <= X"0";
ROM(168) <= X"0";
ROM(169) <= X"7";
ROM(170) <= X"1";
ROM(171) <= X"4";
ROM(172) <= X"1";
ROM(173) <= X"9";
ROM(174) <= X"0";
ROM(175) <= X"0";
	Read_Enable <=  '0' when(CS_L='0' and R_W = '1') else '1';

	
	--process (Clock, Read_Enable, Addr) --Further removed clock signals throughout this process
	process (Read_Enable, Addr)	
	begin  	
		--if(Clock='0') then
			if(Read_Enable = '0') then
			  Data  <= ROM(conv_integer(Addr)); 
		  	else
			  Data <= "ZZZZ";
	      	end if; 
		--else Data <= "ZZZZ";
		--end if;
	
	end process;

	end ROM_176x4_Arch;
